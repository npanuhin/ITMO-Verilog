module Cache (
  input CLK,
  inout wire A1,
  inout wire D1,
  inout wire C1,
  inout wire A2,
  inout wire D2,
  inout wire C2,
  input RESET
);
  always @(RESET) begin

  end
endmodule
