int cache_hits = 0;
int cache_misses = 0;
