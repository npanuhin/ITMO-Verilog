module Hello_World;
  initial begin
    $display("Hello world!");
  end
endmodule
